module (
  input logic in,
  output logic out
);
  
